LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMMAND_DECODER IS
PORT(IR1,IR2:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	EN:IN STD_LOGIC;
	MOVA,MOVB,MOVC,ADD,SUB,OR0,NOT0,RSR,RSL,JMP,JZ,JC,IN0,OUT0,NOP,HALT:OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE structural OF COMMAND_DECODER IS
 SIGNAL temp:STD_LOGIC_VECTOR(15 DOWNTO 0):="0000000000000000";
 SIGNAL prev:STD_LOGIC_VECTOR(3 DOWNTO 0);
 SIGNAL R1,R2:STD_LOGIC_vECTOR(1 DOWNTO 0);
 
BEGIN
 PROCESS(IR1,IR2,EN,temp,prev,R1,R2)
BEGIN
 temp<="0000000000000000";
 prev<=IR1;
 R1<=IR2(3)&IR2(2);
 R2<=IR2(1)&IR2(0);
 
 IF EN='1' THEN
	IF prev="1111" THEN
		IF R1/="11" AND R2/="11" THEN temp<="1000000000000000";
			ELSIF R1="11" AND R2/="11" THEN temp<="0100000000000000";
			ELSIF R1/="11" AND R2="11" THEN temp<="0010000000000000";
		END IF;
		ELSIF prev="1001" THEN temp<="0001000000000000";
		ELSIF prev="0110" THEN temp<="0000100000000000";
		ELSIF prev="1011" THEN temp<="0000010000000000";
		ELSIF prev="0101" THEN temp<="0000001000000000";
		ELSIF prev="1010" THEN
			IF R2="00" THEN temp<=	 "0000000100000000";
			ELSIF R2="11" THEN temp<="0000000010000000";
			END IF;
		ELSIF prev="0011" THEN
			IF (R1="00" AND R2="00") THEN temp<="0000000001000000";
			ELSIF (R1="00" AND R2="01") THEN temp<="0000000000100000";
			ELSIF (R1="00" AND R2="10") THEN temp<="0000000000010000";
			END IF;
		ELSIF prev="0010" THEN temp<="0000000000001000";
		ELSIF prev="0100" THEN temp<="0000000000000100";
		ELSIF (prev="0111" AND R1="00" AND R2="00") THEN temp<="0000000000000010";
		ELSIF (prev="1000" AND R1="00" AND R2="00") THEN temp<="0000000000000001";
		END IF;
	END IF;
		IF temp(15)='1' THEN MOVA<='1';
		ELSE MOVA<='0';
		END IF;
		IF temp(14)='1' THEN MOVB<='1';
		ELSE MOVB<='0';
		END IF;
		IF temp(13)='1' THEN MOVC<='1';
		ELSE MOVC<='0';
		END IF;
		IF temp(12)='1'  THEN ADD<='1';
		ELSE ADD<='0';
		END IF;
		IF temp(11)='1'  THEN SUB<='1';
		ELSE SUB<='0';
		END IF;
		IF temp(10)='1'  THEN OR0<='1';
		ELSE OR0<='0';
		END IF;
		IF temp(9)='1'  THEN NOT0<='1';
		ELSE NOT0<='0';
		END IF;
		IF temp(8)='1'  THEN RSR<='1';
		ELSE RSR<='0';
		END IF;
		IF temp(7)='1'  THEN RSL<='1';
		ELSE RSL<='0';
		END IF;
		IF temp(6)='1'  THEN JMP<='1';
		ELSE JMP<='0';
		END IF;
		IF temp(5)='1'  THEN JZ<='1';
		ELSE JZ<='0';
		END IF;
		IF temp(4)='1'  THEN JC<='1';
		ELSE JC<='0';
		END IF;
		IF temp(3)='1'  THEN IN0<='1';
		ELSE IN0<='0';
		END IF;
		IF temp(2)='1'  THEN OUT0<='1';
		ELSE OUT0<='0';
		END IF;
		IF temp(1)='1'  THEN NOP<='1';
		ELSE NOP<='0';
		END IF;
		IF temp(0)='1'  THEN HALT<='1';
		ELSE HALT<='0';
		END IF;
	END PROCESS;
END structural;